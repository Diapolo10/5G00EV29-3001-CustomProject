.title KiCad schematic
C2 GND Net-_C2-Pad2_ C
C1 GND Net-_C1-Pad2_ C
BT1 Net-_BT1-Pad1_ GND Battery
R1 NC_01 NC_02 10k resistor
SW1 Net-_SW1-Pad1_ Net-_BT1-Pad1_ Reset
U1 Net-_SW1-Pad1_ NC_03 NC_04 NC_05 NC_06 NC_07 Net-_BT1-Pad1_ GND Net-_C1-Pad2_ Net-_C2-Pad2_ NC_08 NC_09 NC_10 NC_11 NC_12 NC_13 NC_14 NC_15 NC_16 NC_17 NC_18 GND NC_19 NC_20 NC_21 NC_22 NC_23 NC_24 ATmega328P-PU
Y1 Net-_C1-Pad2_ Net-_C2-Pad2_ Crystal
.end
